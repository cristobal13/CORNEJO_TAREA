

module ALU 
(
	input [3:0] ALUOperation,
	input [31:0] A,
	input [31:0] B,
	input [4:0] shamt,
	output reg Zero,
	output reg [31:0]ALUResult
);

localparam AND = 4'b0000;
localparam OR  = 4'b0001;
localparam NOR = 4'b0010;
localparam ADD = 4'b0011;
localparam SUB = 4'b0100;
localparam SLL = 4'b0110;
localparam SRL = 4'b0111;



   
   always @ (A or B or ALUOperation)
     begin
		case (ALUOperation)
		
		  ADD: // add
			ALUResult= A + B;
		  SUB: // sub
			ALUResult=A - B;
		   AND: //add
			ALUResult = A & B;
			OR://or
			ALUResult= A | B;
			NOR://nor
			ALUResult= ~(A|B);
			SLL:
			ALUResult= B<< shamt;
			SRL:
			ALUResult= B>> shamt;
			
			
			
			
			

		default:
			ALUResult= 0;
		endcase // case(control)
		Zero = (ALUResult==0) ? 1'b1 : 1'b0;
     end // always @ (A or B or control)
endmodule // ALU